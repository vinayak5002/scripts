// module dff(input j, input k, input clk, output q)